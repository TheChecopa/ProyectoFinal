module branch
(
	input zero, pcsrc,
	output salida
	
);

assign salida = zero & pcsrc;


endmodule 